// File Name: regfile_assign.sv
// Engineer:  Tarun Prakash
// Description:  Code used in regfile.sv for assignment
//          
///////////////////////////////////////////////////////////////////

config_bits[OPBIAS1] <= 8'h00; 
config_bits[OPBIAS2] <= 8'h00;
config_bits[S_PIXEL_EN] <= 8'h00;
config_bits[S_PIXEL_ROW] <= 8'h00;
config_bits[S_PIXEL_COL] <= 8'h00;
config_bits[PIXEL_DISABLE] <= 8'h01;
config_bits[CDS]   <= 8'h00;
config_bits[REG8]  <= 8'h00;      
config_bits[REG9]  <= 8'h00;      
config_bits[REG10] <= 8'h00;      
config_bits[REG11] <= 8'h00;      
config_bits[REG12] <= 8'h02;      //spare0
config_bits[REG13] <= 8'h09;      //spare1
config_bits[REG14] <= 8'h00;      
config_bits[REG15] <= 8'h00;      
config_bits[REG16] <= 8'h00;      

